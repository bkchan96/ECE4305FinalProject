`timescale 1ns / 1ps

module symbol
    (
        input [2:0] value,
        input [9:0] pixel_x, pixel_y,
        input [9:0] top_left_x, top_left_y,
        output on,
        output reg [11:0] color
    );
    
    // load in and declare position and sizing of number
    localparam FOOTPRINT = 32;                                 
    wire [9:0] C_X_L = top_left_x;                   
    wire [9:0] C_Y_T = top_left_y;                  
    wire [9:0] C_X_R = C_X_L + FOOTPRINT - 1;
    wire [9:0] C_Y_B = C_Y_T + FOOTPRINT - 1;
    
    // declare signals to check
    wire [4:0] rom_addr, rom_col;
    wire rom_bit;
    wire sq_on;
    reg [0:31] rom_data;
    
    // check current position of pixel
    assign rom_addr = pixel_y[4:0] - C_Y_T[4:0];
    assign rom_col = pixel_x[4:0] - C_X_L[4:0];
    assign rom_bit = rom_data[rom_col];
    
    // enable on if within foot print
    assign sq_on =
       (C_X_L<=pixel_x) && (pixel_x<=C_X_R) &&
       (C_Y_T<=pixel_y) && (pixel_y<=C_Y_B);
    
    //enable
    assign on = sq_on & rom_bit;
    
    // determine number to output
    always @* begin
        if (value == 0) begin
            color = 12'b111100000000; // red
            case (rom_addr)
                5'd0:  rom_data <=    32'b0000000000000000_0000000000000000;
                5'd1:  rom_data <=    32'b0000000000000000_0000000000000000;
                5'd2:  rom_data <=    32'b0000000000000000_0000000000000000;
                5'd3:  rom_data <=    32'b0000000000000000_0000000000000000;
                5'd4:  rom_data <=    32'b0000111111111111_1111111111110000;
                5'd5:  rom_data <=    32'b0000111111111111_1111111111110000;
                5'd6:  rom_data <=    32'b0000111111111111_1111111111110000;
                5'd7:  rom_data <=    32'b0000111111111111_1111111111110000;
                5'd8:  rom_data <=    32'b0000111111111111_1111111111110000;
                5'd9:  rom_data <=    32'b0000111111111111_1111111111110000;
                5'd10: rom_data <=    32'b0000111111111111_1111111111110000;
                5'd11: rom_data <=    32'b0000111111111111_1111111111110000;
                5'd12: rom_data <=    32'b0000111111111111_1111111111110000;
                5'd13: rom_data <=    32'b0000111111111111_1111111111110000;
                5'd14: rom_data <=    32'b0000111111111111_1111111111110000;         
                5'd15: rom_data <=    32'b0000111111111111_1111111111110000;
                5'd16: rom_data <=    32'b0000111111111111_1111111111110000;   
                5'd17: rom_data <=    32'b0000111111111111_1111111111110000;   
                5'd18: rom_data <=    32'b0000111111111111_1111111111110000;   
                5'd19: rom_data <=    32'b0000111111111111_1111111111110000;   
                5'd20: rom_data <=    32'b0000111111111111_1111111111110000;   
                5'd21: rom_data <=    32'b0000111111111111_1111111111110000;   
                5'd22: rom_data <=    32'b0000111111111111_1111111111110000;   
                5'd23: rom_data <=    32'b0000111111111111_1111111111110000;   
                5'd24: rom_data <=    32'b0000111111111111_1111111111110000;
                5'd25: rom_data <=    32'b0000111111111111_1111111111110000;   
                5'd26: rom_data <=    32'b0000111111111111_1111111111110000;   
                5'd27: rom_data <=    32'b0000111111111111_1111111111110000;   
                5'd28: rom_data <=    32'b0000000000000000_0000000000000000;   
                5'd29: rom_data <=    32'b0000000000000000_0000000000000000;
                5'd30: rom_data <=    32'b0000000000000000_0000000000000000;
                5'd31: rom_data <=    32'b0000000000000000_0000000000000000;
            endcase
        end
        else if (value == 1) begin
            color = 12'b111111110000; // yellow
            case (rom_addr)
                5'd0:  rom_data <=    32'b0000000000000000_0000000000000000;
                5'd1:  rom_data <=    32'b0000000000000000_0000000000000000;
                5'd2:  rom_data <=    32'b0000000000000001_1000000000000000;
                5'd3:  rom_data <=    32'b0000000000000011_1100000000000000;
                5'd4:  rom_data <=    32'b0000000000000111_1110000000000000;
                5'd5:  rom_data <=    32'b0000000000001111_1111000000000000;
                5'd6:  rom_data <=    32'b0000000000011111_1111100000000000;
                5'd7:  rom_data <=    32'b0000000000111111_1111110000000000;
                5'd8:  rom_data <=    32'b0000000001111111_1111111000000000;
                5'd9:  rom_data <=    32'b0000000011111111_1111111100000000;
                5'd10: rom_data <=    32'b0000000111111111_1111111110000000;
                5'd11: rom_data <=    32'b0000001111111111_1111111111000000;
                5'd12: rom_data <=    32'b0000011111111111_1111111111100000;
                5'd13: rom_data <=    32'b0000111111111111_1111111111110000;
                5'd14: rom_data <=    32'b0001111111111111_1111111111111000;         
                5'd15: rom_data <=    32'b0011111111111111_1111111111111100;
                5'd16: rom_data <=    32'b0011111111111111_1111111111111100;   
                5'd17: rom_data <=    32'b0001111111111111_1111111111111000;   
                5'd18: rom_data <=    32'b0000111111111111_1111111111110000;   
                5'd19: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd20: rom_data <=    32'b0000001111111111_1111111111000000;   
                5'd21: rom_data <=    32'b0000000111111111_1111111110000000;   
                5'd22: rom_data <=    32'b0000000011111111_1111111100000000;   
                5'd23: rom_data <=    32'b0000000001111111_1111111000000000;   
                5'd24: rom_data <=    32'b0000000000111111_1111110000000000;
                5'd25: rom_data <=    32'b0000000000011111_1111100000000000;   
                5'd26: rom_data <=    32'b0000000000001111_1111000000000000;   
                5'd27: rom_data <=    32'b0000000000000111_1110000000000000;   
                5'd28: rom_data <=    32'b0000000000000011_1100000000000000;   
                5'd29: rom_data <=    32'b0000000000000001_1000000000000000;
                5'd30: rom_data <=    32'b0000000000000000_0000000000000000;
                5'd31: rom_data <=    32'b0000000000000000_0000000000000000;
            endcase
        end
        else if (value == 2) begin
            color = 12'b000000001111; // blue
            case (rom_addr)
                5'd0:  rom_data <=    32'b0000000000000000_0000000000000000;
                5'd1:  rom_data <=    32'b0000000000000000_0000000000000000;
                5'd2:  rom_data <=    32'b0000000000000001_1000000000000000;
                5'd3:  rom_data <=    32'b0000000000000011_1100000000000000;
                5'd4:  rom_data <=    32'b0000011111111111_1111111111100000;
                5'd5:  rom_data <=    32'b0000011111111111_1111111111100000;
                5'd6:  rom_data <=    32'b0000011111111111_1111111111100000;
                5'd7:  rom_data <=    32'b0000011111111111_1111111111100000;
                5'd8:  rom_data <=    32'b0000011111111111_1111111111100000;
                5'd9:  rom_data <=    32'b0000011111111111_1111111111100000;
                5'd10: rom_data <=    32'b0000011111111111_1111111111100000;
                5'd11: rom_data <=    32'b0000011111111111_1111111111100000;
                5'd12: rom_data <=    32'b0000011111111111_1111111111100000;
                5'd13: rom_data <=    32'b0000111111111111_1111111111100000;
                5'd14: rom_data <=    32'b0001111111111111_1111111111110000;         
                5'd15: rom_data <=    32'b0011111111111111_1111111111111000;
                5'd16: rom_data <=    32'b0011111111111111_1111111111111100;   
                5'd17: rom_data <=    32'b0001111111111111_1111111111111000;   
                5'd18: rom_data <=    32'b0000111111111111_1111111111110000;   
                5'd19: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd20: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd21: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd22: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd23: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd24: rom_data <=    32'b0000011111111111_1111111111100000;
                5'd25: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd26: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd27: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd28: rom_data <=    32'b0000000000000011_1100000000000000;   
                5'd29: rom_data <=    32'b0000000000000001_1000000000000000;
                5'd30: rom_data <=    32'b0000000000000000_0000000000000000;
                5'd31: rom_data <=    32'b0000000000000000_0000000000000000;
            endcase
        end
        else if (value == 3) begin
            color = 12'b000000010000; // green
            case (rom_addr)
                5'd0:  rom_data <=    32'b0000000000000000_0000000000000000;
                5'd1:  rom_data <=    32'b0000000000000000_0000000000000000;
                5'd2:  rom_data <=    32'b0000000000000001_1000000000000000;
                5'd3:  rom_data <=    32'b0000000000000011_1100000000000000;
                5'd4:  rom_data <=    32'b0000011111111111_1111111111100000;
                5'd5:  rom_data <=    32'b0000011111111111_1111111111100000;
                5'd6:  rom_data <=    32'b0000011111111111_1111111111100000;
                5'd7:  rom_data <=    32'b0000011111111111_1111111111100000;
                5'd8:  rom_data <=    32'b0000011111111111_1111111111100000;
                5'd9:  rom_data <=    32'b0000011111111111_1111111111100000;
                5'd10: rom_data <=    32'b0000011111111111_1111111111100000;
                5'd11: rom_data <=    32'b0000011111111111_1111111111100000;
                5'd12: rom_data <=    32'b0000011111111111_1111111111100000;
                5'd13: rom_data <=    32'b0000111111111111_1111111111100000;
                5'd14: rom_data <=    32'b0001111111111111_1111111111110000;         
                5'd15: rom_data <=    32'b0011111111111111_1111111111111000;
                5'd16: rom_data <=    32'b0011111111111111_1111111111111100;   
                5'd17: rom_data <=    32'b0001111111111111_1111111111111000;   
                5'd18: rom_data <=    32'b0000111111111111_1111111111110000;   
                5'd19: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd20: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd21: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd22: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd23: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd24: rom_data <=    32'b0000011111111111_1111111111100000;
                5'd25: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd26: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd27: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd28: rom_data <=    32'b0000000000000011_1100000000000000;   
                5'd29: rom_data <=    32'b0000000000000001_1000000000000000;
                5'd30: rom_data <=    32'b0000000000000000_0000000000000000;
                5'd31: rom_data <=    32'b0000000000000000_0000000000000000;
            endcase
        end
        else if (value == 4) begin
            color = 12'b000000000000; // black
            case (rom_addr)
                5'd0:  rom_data <=    32'b0000000000000000_0000000000000000;
                5'd1:  rom_data <=    32'b0000000000000000_0000000000000000;
                5'd2:  rom_data <=    32'b0000000000000001_1000000000000000;
                5'd3:  rom_data <=    32'b0000000000000011_1100000000000000;
                5'd4:  rom_data <=    32'b0000000000000111_1110000000000000;
                5'd5:  rom_data <=    32'b0000000000001111_1111000000000000;
                5'd6:  rom_data <=    32'b0000000000011111_1111100000000000;
                5'd7:  rom_data <=    32'b0000000000111111_1111110000000000;
                5'd8:  rom_data <=    32'b0000000001111111_1111111000000000;
                5'd9:  rom_data <=    32'b0000000011111111_1111111100000000;
                5'd10: rom_data <=    32'b0000000111111111_1111111110000000;
                5'd11: rom_data <=    32'b0000001111111111_1111111111000000;
                5'd12: rom_data <=    32'b0000011111111111_1111111111100000;
                5'd13: rom_data <=    32'b0000111111111111_1111111111110000;
                5'd14: rom_data <=    32'b0001111111111111_1111111111111000;         
                5'd15: rom_data <=    32'b0011111111111111_1111111111111100;
                5'd16: rom_data <=    32'b0011111111111111_1111111111111100;   
                5'd17: rom_data <=    32'b0001111111111111_1111111111111000;   
                5'd18: rom_data <=    32'b0000111111111111_1111111111110000;   
                5'd19: rom_data <=    32'b0000011111111111_1111111111100000;   
                5'd20: rom_data <=    32'b0000001111111111_1111111111000000;   
                5'd21: rom_data <=    32'b0000000111111111_1111111110000000;   
                5'd22: rom_data <=    32'b0000000011111111_1111111100000000;   
                5'd23: rom_data <=    32'b0000000001111111_1111111000000000;   
                5'd24: rom_data <=    32'b0000000000111111_1111110000000000;
                5'd25: rom_data <=    32'b0000000000011111_1111100000000000;   
                5'd26: rom_data <=    32'b0000000000001111_1111000000000000;   
                5'd27: rom_data <=    32'b0000000000000111_1110000000000000;   
                5'd28: rom_data <=    32'b0000000000000011_1100000000000000;   
                5'd29: rom_data <=    32'b0000000000000001_1000000000000000;
                5'd30: rom_data <=    32'b0000000000000000_0000000000000000;
                5'd31: rom_data <=    32'b0000000000000000_0000000000000000;
            endcase
        end
        // test case for empty
        else if (value == 7) begin
            color = 12'b111111111111; // white
            case (rom_addr)
                5'd0:  rom_data <=    32'b1111111111111111_1111111111111111;
                5'd1:  rom_data <=    32'b1111111111111111_1111111111111111;
                5'd2:  rom_data <=    32'b1111111111111111_1111111111111111;
                5'd3:  rom_data <=    32'b1111111111111111_1111111111111111;
                5'd4:  rom_data <=    32'b1111111111111111_1111111111111111;
                5'd5:  rom_data <=    32'b1111111111111111_1111111111111111;
                5'd6:  rom_data <=    32'b1111111111111111_1111111111111111;
                5'd7:  rom_data <=    32'b1111111111111111_1111111111111111;
                5'd8:  rom_data <=    32'b1111111111111111_1111111111111111;
                5'd9:  rom_data <=    32'b1111111111111111_1111111111111111;
                5'd10: rom_data <=    32'b1111111111111111_1111111111111111;
                5'd11: rom_data <=    32'b1111111111111111_1111111111111111;
                5'd12: rom_data <=    32'b1111111111111111_1111111111111111;
                5'd13: rom_data <=    32'b1111111111111111_1111111111111111;
                5'd14: rom_data <=    32'b1111111111111111_1111111111111111;         
                5'd15: rom_data <=    32'b1111111111111111_1111111111111111;
                5'd16: rom_data <=    32'b1111111111111111_1111111111111111;   
                5'd17: rom_data <=    32'b1111111111111111_1111111111111111;   
                5'd18: rom_data <=    32'b1111111111111111_1111111111111111;   
                5'd19: rom_data <=    32'b1111111111111111_1111111111111111;   
                5'd20: rom_data <=    32'b1111111111111111_1111111111111111;   
                5'd21: rom_data <=    32'b1111111111111111_1111111111111111;   
                5'd22: rom_data <=    32'b1111111111111111_1111111111111111;   
                5'd23: rom_data <=    32'b1111111111111111_1111111111111111;   
                5'd24: rom_data <=    32'b1111111111111111_1111111111111111;
                5'd25: rom_data <=    32'b1111111111111111_1111111111111111;   
                5'd26: rom_data <=    32'b1111111111111111_1111111111111111;   
                5'd27: rom_data <=    32'b1111111111111111_1111111111111111;   
                5'd28: rom_data <=    32'b1111111111111111_1111111111111111;   
                5'd29: rom_data <=    32'b1111111111111111_1111111111111111;
                5'd30: rom_data <=    32'b1111111111111111_1111111111111111;
                5'd31: rom_data <=    32'b1111111111111111_1111111111111111;
            endcase
        end
    end
endmodule